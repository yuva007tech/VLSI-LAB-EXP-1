module full_subtractor(a, b, c,D, Bout);

input a, b, c;

output D, Bout;

assign D = a^b^c;

assign Bout = (~a & b) | (~(a^ b) & c);

endmodule
